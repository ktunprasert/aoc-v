module aoc2024_day1

const input_file = '1.txt'
const example_file = '1e.txt'

fn parse_input() {}
